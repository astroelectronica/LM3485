.title KiCad schematic
.include "C:/AE/LM3485/_models/6TPC100M.lib"
.include "C:/AE/LM3485/_models/ASLL_865060543003_22uF.lib"
.include "C:/AE/LM3485/_models/C2012C0G2A102J060AA_p.mod"
.include "C:/AE/LM3485/_models/C2012X7R2A104K125AA_p.mod"
.include "C:/AE/LM3485/_models/CGJ4C2C0G2A101J060AA_p.mod"
.include "C:/AE/LM3485/_models/MBRS130T3.LIB"
.include "C:/AE/LM3485/_models/PD_7345_7447773220_22u.lib"
.include "C:/AE/LM3485/_models/ZXMP7A17K.lib"
.include "C:/AE/LM3485/_models/lm3485.lib"
R1 VCC /ADJ {RADJ}
XU2 VCC /ADJ C2012C0G2A102J060AA_p
XU3 VCC 0 C2012X7R2A104K125AA_p
XU4 VCC 0 C2012X7R2A104K125AA_p
R2 /OUT /FB {RFBU}
XU8 /OUT 0 6TPC100M
R3 /FB 0 {RFBB}
I1 /OUT 0 DC {ILOAD} 
XU9 /OUT 0 C2012X7R2A104K125AA_p
XU5 /SENSE 0 /FB /ADJ /G VCC LM3485
D1 0 /SENSE Dmbrs130t3
XU7 /SENSE /OUT PD_7345_7447773220_22u
XU6 /OUT /FB CGJ4C2C0G2A101J060AA_p
XU10 /SENSE /G VCC ZXMP7A17K
XU1 VCC 0 ASLL_865060543003_22uF
V1 VCC 0 DC {VIN} 
.end
